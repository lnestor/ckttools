

module c1908
(
  N1,
  N4,
  N7,
  N10,
  N13,
  N16,
  N19,
  N22,
  N25,
  N28,
  N31,
  N34,
  N37,
  N40,
  N43,
  N46,
  N49,
  N53,
  N56,
  N60,
  N63,
  N66,
  N69,
  N72,
  N76,
  N79,
  N82,
  N85,
  N88,
  N91,
  N94,
  N99,
  N104,
  N2753,
  N2754,
  N2755,
  N2756,
  N2762,
  N2767,
  N2768,
  N2779,
  N2780,
  N2781,
  N2782,
  N2783,
  N2784,
  N2785,
  N2786,
  N2787,
  N2811,
  N2886,
  N2887,
  N2888,
  N2889,
  N2890,
  N2891,
  N2892,
  N2899,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_1_8,
  keyIn_1_9
);

  input N1;input N4;input N7;input N10;input N13;input N16;input N19;input N22;input N25;input N28;input N31;input N34;input N37;input N40;input N43;input N46;input N49;input N53;input N56;input N60;input N63;input N66;input N69;input N72;input N76;input N79;input N82;input N85;input N88;input N91;input N94;input N99;input N104;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_1_8;
  input keyIn_1_9;
  output N2753;output N2754;output N2755;output N2756;output N2762;output N2767;output N2768;output N2779;output N2780;output N2781;output N2782;output N2783;output N2784;output N2785;output N2786;output N2787;output N2811;output N2886;output N2887;output N2888;output N2889;output N2890;output N2891;output N2892;output N2899;
  wire N190;wire N194;wire N197;wire N201;wire N206;wire N209;wire N212;wire N216;wire N220;wire N225;wire N229;wire N232;wire N235;wire N239;wire N243;wire N247;wire N251;wire N252;wire N253;wire N256;wire N257;wire N260;wire N263;wire N266;wire N269;wire N272;wire N275;wire N276;wire N277;wire N280;wire N283;wire N290;wire N297;wire N300;wire N303;wire N306;wire N313;wire N316;wire N319;wire N326;wire N331;wire N338;wire N343;wire N346;wire N349;wire N352;wire N355;wire N358;wire N361;wire N364;wire N367;wire N370;wire N373;wire N376;wire N379;wire N382;wire N385;wire N388;wire N534;wire N535;wire N536;wire N537;wire N538;wire N539;wire N540;wire N541;wire N542;wire N543;wire N544;wire N545;wire N546;wire N547;wire N548;wire N549;wire N550;wire N551;wire N552;wire N553;wire N554;wire N555;wire N556;wire N559;wire N562;wire N565;wire N568;wire N571;wire N574;wire N577;wire N580;wire N583;wire N586;wire N589;wire N592;wire N595;wire N598;wire N601;wire N602;wire N603;wire N608;wire N612;wire N616;wire N619;wire N622;wire N625;wire N628;wire N631;wire N634;wire N637;wire N640;wire N643;wire N646;wire N649;wire N652;wire N655;wire N658;wire N661;wire N664;wire N667;wire N670;wire N673;wire N676;wire N679;wire N682;wire N685;wire N688;wire N691;wire N694;wire N697;wire N700;wire N703;wire N706;wire N709;wire N712;wire N715;wire N718;wire N721;wire N724;wire N727;wire N730;wire N733;wire N736;wire N739;wire N742;wire N745;wire N748;wire N751;wire N886;wire N887;wire N888;wire N889;wire N890;wire N891;wire N892;wire N893;wire N894;wire N895;wire N896;wire N897;wire N898;wire N899;wire N903;wire N907;wire N910;wire N913;wire N914;wire N915;wire N916;wire N917;wire N918;wire N919;wire N920;wire N921;wire N922;wire N923;wire N926;wire N935;wire N938;wire N939;wire N942;wire N943;wire N946;wire N947;wire N950;wire N951;wire N954;wire N955;wire N958;wire N959;wire N962;wire N965;wire N968;wire N969;wire N972;wire N973;wire N976;wire N977;wire N980;wire N981;wire N984;wire N985;wire N988;wire N989;wire N990;wire N991;wire N992;wire N993;wire N994;wire N997;wire N998;wire N1001;wire N1002;wire N1003;wire N1004;wire N1005;wire N1006;wire N1007;wire N1008;wire N1009;wire N1010;wire N1013;wire N1016;wire N1019;wire N1022;wire N1025;wire N1028;wire N1031;wire N1034;wire N1037;wire N1040;wire N1043;wire N1046;wire N1049;wire N1054;wire N1055;wire N1063;wire N1064;wire N1067;wire N1068;wire N1119;wire N1120;wire N1121;wire N1122;wire N1128;wire N1129;wire N1130;wire N1131;wire N1132;wire N1133;wire N1148;wire N1149;wire N1150;wire N1151;wire N1152;wire N1153;wire N1154;wire N1155;wire N1156;wire N1157;wire N1158;wire N1159;wire N1160;wire N1161;wire N1162;wire N1163;wire N1164;wire N1167;wire N1168;wire N1171;wire N1188;wire N1205;wire N1206;wire N1207;wire N1208;wire N1209;wire N1210;wire N1211;wire N1212;wire N1213;wire N1214;wire N1215;wire N1216;wire N1217;wire N1218;wire N1219;wire N1220;wire N1221;wire N1222;wire N1223;wire N1224;wire N1225;wire N1226;wire N1227;wire N1228;wire N1229;wire N1230;wire N1231;wire N1232;wire N1235;wire N1238;wire N1239;wire N1240;wire N1241;wire N1242;wire N1243;wire N1246;wire N1249;wire N1252;wire N1255;wire N1258;wire N1261;wire N1264;wire N1267;wire N1309;wire N1310;wire N1311;wire N1312;wire N1313;wire N1314;wire N1315;wire N1316;wire N1317;wire N1318;wire N1319;wire N1322;wire N1327;wire N1328;wire N1334;wire N1344;wire N1345;wire N1346;wire N1348;wire N1349;wire N1350;wire N1351;wire N1352;wire N1355;wire N1358;wire N1361;wire N1364;wire N1367;wire N1370;wire N1373;wire N1376;wire N1379;wire N1383;wire N1386;wire N1387;wire N1388;wire N1389;wire N1390;wire N1393;wire N1396;wire N1397;wire N1398;wire N1399;wire N1409;wire N1412;wire N1413;wire N1416;wire N1419;wire N1433;wire N1434;wire N1438;wire N1439;wire N1440;wire N1443;wire N1444;wire N1445;wire N1446;wire N1447;wire N1448;wire N1451;wire N1452;wire N1453;wire N1454;wire N1455;wire N1456;wire N1457;wire N1458;wire N1459;wire N1460;wire N1461;wire N1462;wire N1463;wire N1464;wire N1468;wire N1469;wire N1470;wire N1471;wire N1472;wire N1475;wire N1476;wire N1478;wire N1481;wire N1484;wire N1487;wire N1488;wire N1489;wire N1490;wire N1491;wire N1492;wire N1493;wire N1494;wire N1495;wire N1496;wire N1498;wire N1499;wire N1500;wire N1501;wire N1504;wire N1510;wire N1513;wire N1514;wire N1517;wire N1520;wire N1521;wire N1522;wire N1526;wire N1527;wire N1528;wire N1529;wire N1530;wire N1531;wire N1532;wire N1534;wire N1537;wire N1540;wire N1546;wire N1554;wire N1557;wire N1561;wire N1567;wire N1568;wire N1569;wire N1571;wire N1576;wire N1588;wire N1591;wire N1593;wire N1594;wire N1595;wire N1596;wire N1600;wire N1603;wire N1606;wire N1609;wire N1612;wire N1615;wire N1620;wire N1623;wire N1635;wire N1636;wire N1638;wire N1639;wire N1640;wire N1643;wire N1647;wire N1651;wire N1658;wire N1661;wire N1664;wire N1671;wire N1672;wire N1675;wire N1677;wire N1678;wire N1679;wire N1680;wire N1681;wire N1682;wire N1683;wire N1685;wire N1688;wire N1697;wire N1701;wire N1706;wire N1707;wire N1708;wire N1709;wire N1710;wire N1711;wire N1712;wire N1713;wire N1714;wire N1717;wire N1720;wire N1721;wire N1723;wire N1727;wire N1728;wire N1730;wire N1731;wire N1734;wire N1740;wire N1741;wire N1742;wire N1746;wire N1747;wire N1748;wire N1751;wire N1759;wire N1761;wire N1762;wire N1763;wire N1764;wire N1768;wire N1769;wire N1772;wire N1773;wire N1774;wire N1777;wire N1783;wire N1784;wire N1785;wire N1786;wire N1787;wire N1788;wire N1791;wire N1792;wire N1795;wire N1796;wire N1798;wire N1801;wire N1802;wire N1807;wire N1808;wire N1809;wire N1810;wire N1812;wire N1815;wire N1818;wire N1821;wire N1822;wire N1823;wire N1824;wire N1825;wire N1826;wire N1827;wire N1830;wire N1837;wire N1838;wire N1841;wire N1848;wire N1849;wire N1850;wire N1852;wire N1855;wire N1856;wire N1857;wire N1858;wire N1864;wire N1865;wire N1866;wire N1869;wire N1872;wire N1875;wire N1878;wire N1879;wire N1882;wire N1883;wire N1884;wire N1885;wire N1889;wire N1895;wire N1896;wire N1897;wire N1898;wire N1902;wire N1910;wire N1911;wire N1912;wire N1913;wire N1915;wire N1919;wire N1920;wire N1921;wire N1922;wire N1923;wire N1924;wire N1927;wire N1930;wire N1933;wire N1936;wire N1937;wire N1938;wire N1941;wire N1942;wire N1944;wire N1947;wire N1950;wire N1953;wire N1958;wire N1961;wire N1965;wire N1968;wire N1975;wire N1976;wire N1977;wire N1978;wire N1979;wire N1980;wire N1985;wire N1987;wire N1999;wire N2000;wire N2002;wire N2003;wire N2004;wire N2005;wire N2006;wire N2007;wire N2008;wire N2009;wire N2012;wire N2013;wire N2014;wire N2015;wire N2016;wire N2018;wire N2019;wire N2020;wire N2021;wire N2022;wire N2023;wire N2024;wire N2025;wire N2026;wire N2027;wire N2030;wire N2033;wire N2036;wire N2037;wire N2038;wire N2039;wire N2040;wire N2041;wire N2042;wire N2047;wire N2052;wire N2055;wire N2060;wire N2061;wire N2062;wire N2067;wire N2068;wire N2071;wire N2076;wire N2077;wire N2078;wire N2081;wire N2086;wire N2089;wire N2104;wire N2119;wire N2129;wire N2143;wire N2148;wire N2151;wire N2196;wire N2199;wire N2202;wire N2205;wire N2214;wire N2215;wire N2216;wire N2217;wire N2222;wire N2223;wire N2224;wire N2225;wire N2226;wire N2227;wire N2228;wire N2229;wire N2230;wire N2231;wire N2232;wire N2233;wire N2234;wire N2235;wire N2236;wire N2237;wire N2240;wire N2241;wire N2244;wire N2245;wire N2250;wire N2253;wire N2256;wire N2257;wire N2260;wire N2263;wire N2266;wire N2269;wire N2272;wire N2279;wire N2286;wire N2297;wire N2315;wire N2326;wire N2340;wire N2353;wire N2361;wire N2375;wire N2384;wire N2385;wire N2386;wire N2426;wire N2427;wire N2537;wire N2540;wire N2543;wire N2546;wire N2549;wire N2552;wire N2555;wire N2558;wire N2561;wire N2564;wire N2567;wire N2570;wire N2573;wire N2576;wire N2594;wire N2597;wire N2600;wire N2603;wire N2606;wire N2611;wire N2614;wire N2617;wire N2620;wire N2627;wire N2628;wire N2629;wire N2630;wire N2631;wire N2632;wire N2633;wire N2634;wire N2639;wire N2642;wire N2645;wire N2648;wire N2651;wire N2655;wire N2658;wire N2661;wire N2664;wire N2669;wire N2670;wire N2671;wire N2672;wire N2673;wire N2674;wire N2675;wire N2676;wire N2682;wire N2683;wire N2688;wire N2689;wire N2690;wire N2691;wire N2710;wire N2720;wire N2721;wire N2722;wire N2723;wire N2724;wire N2725;wire N2726;wire N2727;wire N2728;wire N2729;wire N2730;wire N2731;wire N2732;wire N2733;wire N2734;wire N2735;wire N2736;wire N2737;wire N2738;wire N2739;wire N2740;wire N2741;wire N2742;wire N2743;wire N2744;wire N2745;wire N2746;wire N2747;wire N2750;wire N2757;wire N2758;wire N2759;wire N2760;wire N2761;wire N2763;wire N2764;wire N2765;wire N2766;wire N2773;wire N2776;wire N2788;wire N2789;wire N2800;wire N2807;wire N2808;wire N2809;wire N2810;wire N2812;wire N2815;wire N2818;wire N2821;wire N2824;wire N2827;wire N2828;wire N2829;wire N2843;wire N2846;wire N2850;wire N2851;wire N2852;wire N2853;wire N2854;wire N2857;wire N2858;wire N2859;wire N2860;wire N2861;wire N2862;wire N2863;wire N2866;wire N2867;wire N2868;wire N2869;wire N2870;wire N2871;wire N2872;wire N2873;wire N2874;wire N2875;wire N2876;wire N2877;wire N2878;wire N2879;wire N2880;wire N2881;wire N2882;wire N2883;wire N2895;wire N2896;wire N2897;wire N2898;
  wire sig_comp_0_0;
  wire sig_comp_0_1;
  wire sig_comp_0_2;
  wire sig_comp_0_3;
  wire sig_comp_0_4;
  wire sig_comp_0_5;
  wire sig_comp_0_6;
  wire sig_comp_0_7;
  wire sig_comp_and_0;
  wire const_comp_xor_0_0;
  wire const_comp_xor_0_1;
  wire const_comp_xor_0_2;
  wire const_comp_xor_0_3;
  wire const_comp_xor_0_4;
  wire const_comp_xor_0_5;
  wire const_comp_xor_0_6;
  wire const_comp_xor_0_7;
  wire const_comp_and_0;
  wire mask_and_0;
  wire signal_from_circuit_0;
  wire mux_control_xor_1_0;
  wire mux_control_xor_1_1;
  wire mux_not_1_0;
  wire mux_and0_1_0;
  wire mux_and1_1_0;
  wire mux_not_1_1;
  wire mux_and0_1_1;
  wire mux_and1_1_1;

  not
  NOT1_1
  (
    N190,
    N1
  );


  not
  NOT1_2
  (
    N194,
    N4
  );


  not
  NOT1_3
  (
    N197,
    N7
  );


  not
  NOT1_4
  (
    N201,
    N10
  );


  not
  NOT1_5
  (
    N206,
    N13
  );


  not
  NOT1_6
  (
    N209,
    N16
  );


  not
  NOT1_7
  (
    N212,
    N19
  );


  not
  NOT1_8
  (
    N216,
    N22
  );


  not
  NOT1_9
  (
    N220,
    N25
  );


  not
  NOT1_10
  (
    N225,
    N28
  );


  not
  NOT1_11
  (
    N229,
    N31
  );


  not
  NOT1_12
  (
    N232,
    N34
  );


  not
  NOT1_13
  (
    N235,
    N37
  );


  not
  NOT1_14
  (
    N239,
    N40
  );


  not
  NOT1_15
  (
    N243,
    N43
  );


  not
  NOT1_16
  (
    N247,
    N46
  );


  nand
  NAND2_17
  (
    N251,
    N63,
    N88
  );


  nand
  NAND2_18
  (
    N252,
    N66,
    N91
  );


  not
  NOT1_19
  (
    N253,
    N72
  );


  not
  NOT1_20
  (
    N256,
    N72
  );


  buf
  BUFF1_21
  (
    N257,
    N69
  );


  buf
  BUFF1_22
  (
    N260,
    N69
  );


  not
  NOT1_23
  (
    N263,
    N76
  );


  not
  NOT1_24
  (
    N266,
    N79
  );


  not
  NOT1_25
  (
    N269,
    N82
  );


  not
  NOT1_26
  (
    N272,
    N85
  );


  not
  NOT1_27
  (
    N275,
    N104
  );


  not
  NOT1_28
  (
    N276,
    N104
  );


  not
  NOT1_29
  (
    N277,
    N88
  );


  not
  NOT1_30
  (
    N280,
    N91
  );


  buf
  BUFF1_31
  (
    N283,
    N94
  );


  not
  NOT1_32
  (
    N290,
    N94
  );


  buf
  BUFF1_33
  (
    N297,
    N94
  );


  not
  NOT1_34
  (
    N300,
    N94
  );


  buf
  BUFF1_35
  (
    N303,
    N99
  );


  not
  NOT1_36
  (
    N306,
    N99
  );


  not
  NOT1_37
  (
    N313,
    N99
  );


  buf
  BUFF1_38
  (
    N316,
    N104
  );


  not
  NOT1_39
  (
    N319,
    N104
  );


  buf
  BUFF1_40
  (
    N326,
    N104
  );


  buf
  BUFF1_41
  (
    N331,
    N104
  );


  not
  NOT1_42
  (
    N338,
    N104
  );


  buf
  BUFF1_43
  (
    N343,
    N1
  );


  buf
  BUFF1_44
  (
    N346,
    N4
  );


  buf
  BUFF1_45
  (
    N349,
    N7
  );


  buf
  BUFF1_46
  (
    N352,
    N10
  );


  buf
  BUFF1_47
  (
    N355,
    N13
  );


  buf
  BUFF1_48
  (
    N358,
    N16
  );


  buf
  BUFF1_49
  (
    N361,
    N19
  );


  buf
  BUFF1_50
  (
    N364,
    N22
  );


  buf
  BUFF1_51
  (
    N367,
    N25
  );


  buf
  BUFF1_52
  (
    N370,
    N28
  );


  buf
  BUFF1_53
  (
    N373,
    N31
  );


  buf
  BUFF1_54
  (
    N376,
    N34
  );


  buf
  BUFF1_55
  (
    N379,
    N37
  );


  buf
  BUFF1_56
  (
    N382,
    N40
  );


  buf
  BUFF1_57
  (
    N385,
    N43
  );


  buf
  BUFF1_58
  (
    N388,
    N46
  );


  not
  NOT1_59
  (
    N534,
    N343
  );


  not
  NOT1_60
  (
    N535,
    N346
  );


  not
  NOT1_61
  (
    N536,
    N349
  );


  not
  NOT1_62
  (
    N537,
    N352
  );


  not
  NOT1_63
  (
    N538,
    N355
  );


  not
  NOT1_64
  (
    N539,
    N358
  );


  not
  NOT1_65
  (
    N540,
    N361
  );


  not
  NOT1_66
  (
    N541,
    N364
  );


  not
  NOT1_67
  (
    N542,
    N367
  );


  not
  NOT1_68
  (
    N543,
    N370
  );


  not
  NOT1_69
  (
    N544,
    N373
  );


  not
  NOT1_70
  (
    N545,
    N376
  );


  not
  NOT1_71
  (
    N546,
    N379
  );


  not
  NOT1_72
  (
    N547,
    N382
  );


  not
  NOT1_73
  (
    N548,
    N385
  );


  not
  NOT1_74
  (
    N549,
    N388
  );


  nand
  NAND2_75
  (
    N550,
    N306,
    N331
  );


  nand
  NAND2_76
  (
    N551,
    N306,
    N331
  );


  nand
  NAND2_77
  (
    N552,
    N306,
    N331
  );


  nand
  NAND2_78
  (
    N553,
    N306,
    N331
  );


  nand
  NAND2_79
  (
    N554,
    N306,
    N331
  );


  nand
  NAND2_80
  (
    N555,
    N306,
    N331
  );


  buf
  BUFF1_81
  (
    N556,
    N190
  );


  buf
  BUFF1_82
  (
    N559,
    N194
  );


  buf
  BUFF1_83
  (
    N562,
    N206
  );


  buf
  BUFF1_84
  (
    N565,
    N209
  );


  buf
  BUFF1_85
  (
    N568,
    N225
  );


  buf
  BUFF1_86
  (
    N571,
    N243
  );


  and
  AND2_87
  (
    N574,
    N63,
    N319
  );


  buf
  BUFF1_88
  (
    N577,
    N220
  );


  buf
  BUFF1_89
  (
    N580,
    N229
  );


  buf
  BUFF1_90
  (
    N583,
    N232
  );


  and
  AND2_91
  (
    N586,
    N66,
    N319
  );


  buf
  BUFF1_92
  (
    N589,
    N239
  );


  and
  AND3_93
  (
    N592,
    N49,
    N253,
    N319
  );


  buf
  BUFF1_94
  (
    N595,
    N247
  );


  buf
  BUFF1_95
  (
    N598,
    N239
  );


  nand
  NAND2_96
  (
    N601,
    N326,
    N277
  );


  nand
  NAND2_97
  (
    N602,
    N326,
    N280
  );


  nand
  NAND2_98
  (
    N603,
    N260,
    N72
  );


  nand
  NAND2_99
  (
    N608,
    N260,
    N300
  );


  nand
  NAND2_100
  (
    N612,
    N256,
    N300
  );


  buf
  BUFF1_101
  (
    N616,
    N201
  );


  buf
  BUFF1_102
  (
    N619,
    N216
  );


  buf
  BUFF1_103
  (
    N622,
    N220
  );


  buf
  BUFF1_104
  (
    N625,
    N239
  );


  buf
  BUFF1_105
  (
    N628,
    N190
  );


  buf
  BUFF1_106
  (
    N631,
    N190
  );


  buf
  BUFF1_107
  (
    N634,
    N194
  );


  buf
  BUFF1_108
  (
    N637,
    N229
  );


  buf
  BUFF1_109
  (
    N640,
    N197
  );


  and
  AND3_110
  (
    N643,
    N56,
    N257,
    N319
  );


  buf
  BUFF1_111
  (
    N646,
    N232
  );


  buf
  BUFF1_112
  (
    N649,
    N201
  );


  buf
  BUFF1_113
  (
    N652,
    N235
  );


  and
  AND3_114
  (
    N655,
    N60,
    N257,
    N319
  );


  buf
  BUFF1_115
  (
    N658,
    N263
  );


  buf
  BUFF1_116
  (
    N661,
    N263
  );


  buf
  BUFF1_117
  (
    N664,
    N266
  );


  buf
  BUFF1_118
  (
    N667,
    N266
  );


  buf
  BUFF1_119
  (
    N670,
    N269
  );


  buf
  BUFF1_120
  (
    N673,
    N269
  );


  buf
  BUFF1_121
  (
    N676,
    N272
  );


  buf
  BUFF1_122
  (
    N679,
    N272
  );


  and
  AND2_123
  (
    N682,
    N251,
    N316
  );


  and
  AND2_124
  (
    N685,
    N252,
    N316
  );


  buf
  BUFF1_125
  (
    N688,
    N197
  );


  buf
  BUFF1_126
  (
    N691,
    N197
  );


  buf
  BUFF1_127
  (
    N694,
    N212
  );


  buf
  BUFF1_128
  (
    N697,
    N212
  );


  buf
  BUFF1_129
  (
    N700,
    N247
  );


  buf
  BUFF1_130
  (
    N703,
    N247
  );


  buf
  BUFF1_131
  (
    N706,
    N235
  );


  buf
  BUFF1_132
  (
    N709,
    N235
  );


  buf
  BUFF1_133
  (
    N712,
    N201
  );


  buf
  BUFF1_134
  (
    N715,
    N201
  );


  buf
  BUFF1_135
  (
    N718,
    N206
  );


  buf
  BUFF1_136
  (
    N721,
    N216
  );


  and
  AND3_137
  (
    N724,
    N53,
    N253,
    N319
  );


  buf
  BUFF1_138
  (
    N727,
    N243
  );


  buf
  BUFF1_139
  (
    N730,
    N220
  );


  buf
  BUFF1_140
  (
    N733,
    N220
  );


  buf
  BUFF1_141
  (
    N736,
    N209
  );


  buf
  BUFF1_142
  (
    N739,
    N216
  );


  buf
  BUFF1_143
  (
    N742,
    N225
  );


  buf
  BUFF1_144
  (
    N745,
    N243
  );


  buf
  BUFF1_145
  (
    N748,
    N212
  );


  buf
  BUFF1_146
  (
    N751,
    N225
  );


  not
  NOT1_147
  (
    N886,
    N682
  );


  not
  NOT1_148
  (
    N887,
    N685
  );


  not
  NOT1_149
  (
    N888,
    N616
  );


  not
  NOT1_150
  (
    N889,
    N619
  );


  not
  NOT1_151
  (
    N890,
    N622
  );


  not
  NOT1_152
  (
    N891,
    N625
  );


  not
  NOT1_153
  (
    N892,
    N631
  );


  not
  NOT1_154
  (
    N893,
    N643
  );


  not
  NOT1_155
  (
    N894,
    N649
  );


  not
  NOT1_156
  (
    N895,
    N652
  );


  not
  NOT1_157
  (
    N896,
    N655
  );


  and
  AND2_158
  (
    N897,
    N49,
    N612
  );


  and
  AND2_159
  (
    N898,
    N56,
    N608
  );


  nand
  NAND2_160
  (
    N899,
    N53,
    N612
  );


  nand
  NAND2_161
  (
    N903,
    N60,
    N608
  );


  nand
  NAND2_162
  (
    N907,
    N49,
    N612
  );


  nand
  NAND2_163
  (
    N910,
    N56,
    N608
  );


  not
  NOT1_164
  (
    N913,
    N661
  );


  not
  NOT1_165
  (
    N914,
    N658
  );


  not
  NOT1_166
  (
    N915,
    N667
  );


  not
  NOT1_167
  (
    N916,
    N664
  );


  not
  NOT1_168
  (
    N917,
    N673
  );


  not
  NOT1_169
  (
    N918,
    N670
  );


  not
  NOT1_170
  (
    N919,
    N679
  );


  not
  NOT1_171
  (
    N920,
    N676
  );


  nand
  NAND4_172
  (
    N921,
    N277,
    N297,
    N326,
    N603
  );


  nand
  NAND4_173
  (
    N922,
    N280,
    N297,
    N326,
    N603
  );


  nand
  NAND3_174
  (
    N923,
    N303,
    N338,
    N603
  );


  and
  AND3_175
  (
    N926,
    N303,
    N338,
    N603
  );


  buf
  BUFF1_176
  (
    N935,
    N556
  );


  not
  NOT1_177
  (
    N938,
    N688
  );


  buf
  BUFF1_178
  (
    N939,
    N556
  );


  not
  NOT1_179
  (
    N942,
    N691
  );


  buf
  BUFF1_180
  (
    N943,
    N562
  );


  not
  NOT1_181
  (
    N946,
    N694
  );


  buf
  BUFF1_182
  (
    N947,
    N562
  );


  not
  NOT1_183
  (
    N950,
    N697
  );


  buf
  BUFF1_184
  (
    N951,
    N568
  );


  not
  NOT1_185
  (
    N954,
    N700
  );


  buf
  BUFF1_186
  (
    N955,
    N568
  );


  not
  NOT1_187
  (
    N958,
    N703
  );


  buf
  BUFF1_188
  (
    N959,
    N574
  );


  buf
  BUFF1_189
  (
    N962,
    N574
  );


  buf
  BUFF1_190
  (
    N965,
    N580
  );


  not
  NOT1_191
  (
    N968,
    N706
  );


  buf
  BUFF1_192
  (
    N969,
    N580
  );


  not
  NOT1_193
  (
    N972,
    N709
  );


  buf
  BUFF1_194
  (
    N973,
    N586
  );


  not
  NOT1_195
  (
    N976,
    N712
  );


  buf
  BUFF1_196
  (
    N977,
    N586
  );


  not
  NOT1_197
  (
    N980,
    N715
  );


  buf
  BUFF1_198
  (
    N981,
    N592
  );


  not
  NOT1_199
  (
    N984,
    N628
  );


  buf
  BUFF1_200
  (
    N985,
    N592
  );


  not
  NOT1_201
  (
    N988,
    N718
  );


  not
  NOT1_202
  (
    N989,
    N721
  );


  not
  NOT1_203
  (
    N990,
    N634
  );


  not
  NOT1_204
  (
    N991,
    N724
  );


  not
  NOT1_205
  (
    N992,
    N727
  );


  not
  NOT1_206
  (
    N993,
    N637
  );


  buf
  BUFF1_207
  (
    N994,
    N595
  );


  not
  NOT1_208
  (
    N997,
    N730
  );


  buf
  BUFF1_209
  (
    N998,
    N595
  );


  not
  NOT1_210
  (
    N1001,
    N733
  );


  not
  NOT1_211
  (
    N1002,
    N736
  );


  not
  NOT1_212
  (
    N1003,
    N739
  );


  not
  NOT1_213
  (
    N1004,
    N640
  );


  not
  NOT1_214
  (
    N1005,
    N742
  );


  not
  NOT1_215
  (
    N1006,
    N745
  );


  not
  NOT1_216
  (
    N1007,
    N646
  );


  not
  NOT1_217
  (
    N1008,
    N748
  );


  not
  NOT1_218
  (
    N1009,
    N751
  );


  buf
  BUFF1_219
  (
    N1010,
    N559
  );


  buf
  BUFF1_220
  (
    N1013,
    N559
  );


  buf
  BUFF1_221
  (
    N1016,
    N565
  );


  buf
  BUFF1_222
  (
    N1019,
    N565
  );


  buf
  BUFF1_223
  (
    N1022,
    N571
  );


  buf
  BUFF1_224
  (
    N1025,
    N571
  );


  buf
  BUFF1_225
  (
    N1028,
    N577
  );


  buf
  BUFF1_226
  (
    N1031,
    N577
  );


  buf
  BUFF1_227
  (
    N1034,
    N583
  );


  buf
  BUFF1_228
  (
    N1037,
    N583
  );


  buf
  BUFF1_229
  (
    N1040,
    N589
  );


  buf
  BUFF1_230
  (
    N1043,
    N589
  );


  buf
  BUFF1_231
  (
    N1046,
    N598
  );


  buf
  BUFF1_232
  (
    N1049,
    N598
  );


  nand
  NAND2_233
  (
    N1054,
    N619,
    N888
  );


  nand
  NAND2_234
  (
    N1055,
    N616,
    N889
  );


  nand
  NAND2_235
  (
    N1063,
    N625,
    N890
  );


  nand
  NAND2_236
  (
    N1064,
    N622,
    N891
  );


  nand
  NAND2_237
  (
    N1067,
    N655,
    N895
  );


  nand
  NAND2_238
  (
    N1068,
    N652,
    N896
  );


  nand
  NAND2_239
  (
    N1119,
    N721,
    N988
  );


  nand
  NAND2_240
  (
    N1120,
    N718,
    N989
  );


  nand
  NAND2_241
  (
    N1121,
    N727,
    N991
  );


  nand
  NAND2_242
  (
    N1122,
    N724,
    N992
  );


  nand
  NAND2_243
  (
    N1128,
    N739,
    N1002
  );


  nand
  NAND2_244
  (
    N1129,
    N736,
    N1003
  );


  nand
  NAND2_245
  (
    N1130,
    N745,
    N1005
  );


  nand
  NAND2_246
  (
    N1131,
    N742,
    N1006
  );


  nand
  NAND2_247
  (
    N1132,
    N751,
    N1008
  );


  nand
  NAND2_248
  (
    N1133,
    N748,
    N1009
  );


  not
  NOT1_249
  (
    N1148,
    N939
  );


  not
  NOT1_250
  (
    N1149,
    N935
  );


  nand
  NAND2_251
  (
    N1150,
    N1054,
    N1055
  );


  not
  NOT1_252
  (
    N1151,
    N943
  );


  not
  NOT1_253
  (
    N1152,
    N947
  );


  not
  NOT1_254
  (
    N1153,
    N955
  );


  not
  NOT1_255
  (
    N1154,
    N951
  );


  not
  NOT1_256
  (
    N1155,
    N962
  );


  not
  NOT1_257
  (
    N1156,
    N969
  );


  not
  NOT1_258
  (
    N1157,
    N977
  );


  nand
  NAND2_259
  (
    N1158,
    N1063,
    N1064
  );


  not
  NOT1_260
  (
    N1159,
    N985
  );


  nand
  NAND2_261
  (
    N1160,
    N985,
    N892
  );


  not
  NOT1_262
  (
    N1161,
    N998
  );


  nand
  NAND2_263
  (
    N1162,
    N1067,
    N1068
  );


  not
  NOT1_264
  (
    N1163,
    N899
  );


  buf
  BUFF1_265
  (
    N1164,
    N899
  );


  not
  NOT1_266
  (
    N1167,
    N903
  );


  buf
  BUFF1_267
  (
    N1168,
    N903
  );


  nand
  NAND2_268
  (
    N1171,
    N921,
    N923
  );


  nand
  NAND2_269
  (
    N1188,
    N922,
    N923
  );


  not
  NOT1_270
  (
    N1205,
    N1010
  );


  nand
  NAND2_271
  (
    N1206,
    N1010,
    N938
  );


  not
  NOT1_272
  (
    N1207,
    N1013
  );


  nand
  NAND2_273
  (
    N1208,
    N1013,
    N942
  );


  not
  NOT1_274
  (
    N1209,
    N1016
  );


  nand
  NAND2_275
  (
    N1210,
    N1016,
    N946
  );


  not
  NOT1_276
  (
    N1211,
    N1019
  );


  nand
  NAND2_277
  (
    N1212,
    N1019,
    N950
  );


  not
  NOT1_278
  (
    N1213,
    N1022
  );


  nand
  NAND2_279
  (
    N1214,
    N1022,
    N954
  );


  not
  NOT1_280
  (
    N1215,
    N1025
  );


  nand
  NAND2_281
  (
    N1216,
    N1025,
    N958
  );


  not
  NOT1_282
  (
    N1217,
    N1028
  );


  not
  NOT1_283
  (
    N1218,
    N959
  );


  not
  NOT1_284
  (
    N1219,
    N1031
  );


  not
  NOT1_285
  (
    N1220,
    N1034
  );


  nand
  NAND2_286
  (
    N1221,
    N1034,
    N968
  );


  not
  NOT1_287
  (
    N1222,
    N965
  );


  not
  NOT1_288
  (
    N1223,
    N1037
  );


  nand
  NAND2_289
  (
    N1224,
    N1037,
    N972
  );


  not
  NOT1_290
  (
    N1225,
    N1040
  );


  nand
  NAND2_291
  (
    N1226,
    N1040,
    N976
  );


  not
  NOT1_292
  (
    N1227,
    N973
  );


  not
  NOT1_293
  (
    N1228,
    N1043
  );


  nand
  NAND2_294
  (
    N1229,
    N1043,
    N980
  );


  not
  NOT1_295
  (
    N1230,
    N981
  );


  nand
  NAND2_296
  (
    N1231,
    N981,
    N984
  );


  nand
  NAND2_297
  (
    N1232,
    N1119,
    N1120
  );


  nand
  NAND2_298
  (
    N1235,
    N1121,
    N1122
  );


  not
  NOT1_299
  (
    N1238,
    N1046
  );


  nand
  NAND2_300
  (
    N1239,
    N1046,
    N997
  );


  not
  NOT1_301
  (
    N1240,
    N994
  );


  not
  NOT1_302
  (
    N1241,
    N1049
  );


  nand
  NAND2_303
  (
    N1242,
    N1049,
    N1001
  );


  nand
  NAND2_304
  (
    N1243,
    N1128,
    N1129
  );


  nand
  NAND2_305
  (
    N1246,
    N1130,
    N1131
  );


  nand
  NAND2_306
  (
    N1249,
    N1132,
    N1133
  );


  buf
  BUFF1_307
  (
    N1252,
    N907
  );


  buf
  BUFF1_308
  (
    N1255,
    N907
  );


  buf
  BUFF1_309
  (
    N1258,
    N910
  );


  buf
  BUFF1_310
  (
    N1261,
    N910
  );


  not
  NOT1_311
  (
    N1264,
    N1150
  );


  nand
  NAND2_312
  (
    N1267,
    N631,
    N1159
  );


  nand
  NAND2_313
  (
    N1309,
    N688,
    N1205
  );


  nand
  NAND2_314
  (
    N1310,
    N691,
    N1207
  );


  nand
  NAND2_315
  (
    N1311,
    N694,
    N1209
  );


  nand
  NAND2_316
  (
    N1312,
    N697,
    N1211
  );


  nand
  NAND2_317
  (
    N1313,
    N700,
    N1213
  );


  nand
  NAND2_318
  (
    N1314,
    N703,
    N1215
  );


  nand
  NAND2_319
  (
    N1315,
    N706,
    N1220
  );


  nand
  NAND2_320
  (
    N1316,
    N709,
    N1223
  );


  nand
  NAND2_321
  (
    N1317,
    N712,
    N1225
  );


  nand
  NAND2_322
  (
    N1318,
    N715,
    N1228
  );


  not
  NOT1_323
  (
    N1319,
    N1158
  );


  nand
  NAND2_324
  (
    N1322,
    N628,
    N1230
  );


  nand
  NAND2_325
  (
    N1327,
    N730,
    N1238
  );


  nand
  NAND2_326
  (
    N1328,
    N733,
    N1241
  );


  not
  NOT1_327
  (
    N1334,
    N1162
  );


  nand
  NAND2_328
  (
    N1344,
    N1267,
    N1160
  );


  nand
  NAND2_329
  (
    N1345,
    N1249,
    N894
  );


  not
  NOT1_330
  (
    N1346,
    N1249
  );


  not
  NOT1_331
  (
    N1348,
    N1255
  );


  not
  NOT1_332
  (
    N1349,
    N1252
  );


  not
  NOT1_333
  (
    N1350,
    N1261
  );


  not
  NOT1_334
  (
    N1351,
    N1258
  );


  nand
  NAND2_335
  (
    N1352,
    N1309,
    N1206
  );


  nand
  NAND2_336
  (
    N1355,
    N1310,
    N1208
  );


  nand
  NAND2_337
  (
    N1358,
    N1311,
    N1210
  );


  nand
  NAND2_338
  (
    N1361,
    N1312,
    N1212
  );


  nand
  NAND2_339
  (
    N1364,
    N1313,
    N1214
  );


  nand
  NAND2_340
  (
    N1367,
    N1314,
    N1216
  );


  nand
  NAND2_341
  (
    N1370,
    N1315,
    N1221
  );


  nand
  NAND2_342
  (
    N1373,
    N1316,
    N1224
  );


  nand
  NAND2_343
  (
    N1376,
    N1317,
    N1226
  );


  nand
  NAND2_344
  (
    N1379,
    N1318,
    N1229
  );


  nand
  NAND2_345
  (
    N1383,
    N1322,
    N1231
  );


  not
  NOT1_346
  (
    N1386,
    N1232
  );


  nand
  NAND2_347
  (
    N1387,
    N1232,
    N990
  );


  not
  NOT1_348
  (
    N1388,
    N1235
  );


  nand
  NAND2_349
  (
    N1389,
    N1235,
    N993
  );


  nand
  NAND2_350
  (
    N1390,
    N1327,
    N1239
  );


  nand
  NAND2_351
  (
    N1393,
    N1328,
    N1242
  );


  not
  NOT1_352
  (
    N1396,
    N1243
  );


  nand
  NAND2_353
  (
    N1397,
    N1243,
    N1004
  );


  not
  NOT1_354
  (
    N1398,
    N1246
  );


  nand
  NAND2_355
  (
    N1399,
    N1246,
    N1007
  );


  not
  NOT1_356
  (
    N1409,
    N1319
  );


  nand
  NAND2_357
  (
    N1412,
    N649,
    N1346
  );


  not
  NOT1_358
  (
    N1413,
    N1334
  );


  buf
  BUFF1_359
  (
    N1416,
    N1264
  );


  buf
  BUFF1_360
  (
    N1419,
    N1264
  );


  nand
  NAND2_361
  (
    N1433,
    N634,
    N1386
  );


  nand
  NAND2_362
  (
    N1434,
    N637,
    N1388
  );


  nand
  NAND2_363
  (
    N1438,
    N640,
    N1396
  );


  nand
  NAND2_364
  (
    N1439,
    N646,
    N1398
  );


  not
  NOT1_365
  (
    N1440,
    N1344
  );


  nand
  NAND2_366
  (
    N1443,
    N1355,
    N1148
  );


  not
  NOT1_367
  (
    N1444,
    N1355
  );


  nand
  NAND2_368
  (
    N1445,
    N1352,
    N1149
  );


  not
  NOT1_369
  (
    N1446,
    N1352
  );


  nand
  NAND2_370
  (
    N1447,
    N1358,
    N1151
  );


  not
  NOT1_371
  (
    N1448,
    N1358
  );


  nand
  NAND2_372
  (
    N1451,
    N1361,
    N1152
  );


  not
  NOT1_373
  (
    N1452,
    N1361
  );


  nand
  NAND2_374
  (
    N1453,
    N1367,
    N1153
  );


  not
  NOT1_375
  (
    N1454,
    N1367
  );


  nand
  NAND2_376
  (
    N1455,
    N1364,
    N1154
  );


  not
  NOT1_377
  (
    N1456,
    N1364
  );


  nand
  NAND2_378
  (
    N1457,
    N1373,
    N1156
  );


  not
  NOT1_379
  (
    N1458,
    N1373
  );


  nand
  NAND2_380
  (
    N1459,
    N1379,
    N1157
  );


  not
  NOT1_381
  (
    N1460,
    N1379
  );


  not
  NOT1_382
  (
    N1461,
    N1383
  );


  nand
  NAND2_383
  (
    N1462,
    N1393,
    N1161
  );


  not
  NOT1_384
  (
    N1463,
    N1393
  );


  nand
  NAND2_385
  (
    N1464,
    N1345,
    N1412
  );


  not
  NOT1_386
  (
    N1468,
    N1370
  );


  nand
  NAND2_387
  (
    N1469,
    N1370,
    N1222
  );


  not
  NOT1_388
  (
    N1470,
    N1376
  );


  nand
  NAND2_389
  (
    N1471,
    N1376,
    N1227
  );


  nand
  NAND2_390
  (
    N1472,
    N1387,
    N1433
  );


  not
  NOT1_391
  (
    N1475,
    N1390
  );


  nand
  NAND2_392
  (
    N1476,
    N1390,
    N1240
  );


  nand
  NAND2_393
  (
    N1478,
    N1389,
    N1434
  );


  nand
  NAND2_394
  (
    N1481,
    N1399,
    N1439
  );


  nand
  NAND2_395
  (
    N1484,
    N1397,
    N1438
  );


  nand
  NAND2_396
  (
    N1487,
    N939,
    N1444
  );


  nand
  NAND2_397
  (
    N1488,
    N935,
    N1446
  );


  nand
  NAND2_398
  (
    N1489,
    N943,
    N1448
  );


  not
  NOT1_399
  (
    N1490,
    N1419
  );


  not
  NOT1_400
  (
    N1491,
    N1416
  );


  nand
  NAND2_401
  (
    N1492,
    N947,
    N1452
  );


  nand
  NAND2_402
  (
    N1493,
    N955,
    N1454
  );


  nand
  NAND2_403
  (
    N1494,
    N951,
    N1456
  );


  nand
  NAND2_404
  (
    N1495,
    N969,
    N1458
  );


  nand
  NAND2_405
  (
    N1496,
    N977,
    N1460
  );


  nand
  NAND2_406
  (
    N1498,
    N998,
    N1463
  );


  not
  NOT1_407
  (
    N1499,
    N1440
  );


  nand
  NAND2_408
  (
    N1500,
    N965,
    N1468
  );


  nand
  NAND2_409
  (
    N1501,
    N973,
    N1470
  );


  nand
  NAND2_410
  (
    N1504,
    N994,
    N1475
  );


  not
  NOT1_411
  (
    N1510,
    N1464
  );


  nand
  NAND2_412
  (
    N1513,
    N1443,
    N1487
  );


  nand
  NAND2_413
  (
    N1514,
    N1445,
    N1488
  );


  nand
  NAND2_414
  (
    N1517,
    N1447,
    N1489
  );


  nand
  NAND2_415
  (
    N1520,
    N1451,
    N1492
  );


  nand
  NAND2_416
  (
    N1521,
    N1453,
    N1493
  );


  nand
  NAND2_417
  (
    N1522,
    N1455,
    N1494
  );


  nand
  NAND2_418
  (
    N1526,
    N1457,
    N1495
  );


  nand
  NAND2_419
  (
    N1527,
    N1459,
    N1496
  );


  not
  NOT1_420
  (
    N1528,
    N1472
  );


  nand
  NAND2_421
  (
    N1529,
    N1462,
    N1498
  );


  not
  NOT1_422
  (
    N1530,
    N1478
  );


  not
  NOT1_423
  (
    N1531,
    N1481
  );


  not
  NOT1_424
  (
    N1532,
    N1484
  );


  nand
  NAND2_425
  (
    N1534,
    N1471,
    N1501
  );


  nand
  NAND2_426
  (
    N1537,
    N1469,
    N1500
  );


  nand
  NAND2_427
  (
    N1540,
    N1476,
    N1504
  );


  not
  NOT1_428
  (
    N1546,
    N1513
  );


  not
  NOT1_429
  (
    N1554,
    N1521
  );


  not
  NOT1_430
  (
    N1557,
    N1526
  );


  not
  NOT1_431
  (
    N1561,
    N1520
  );


  nand
  NAND2_432
  (
    N1567,
    N1484,
    N1531
  );


  nand
  NAND2_433
  (
    N1568,
    N1481,
    N1532
  );


  not
  NOT1_434
  (
    N1569,
    N1510
  );


  not
  NOT1_435
  (
    N1571,
    N1527
  );


  not
  NOT1_436
  (
    N1576,
    N1529
  );


  buf
  BUFF1_437
  (
    N1588,
    N1522
  );


  not
  NOT1_438
  (
    N1591,
    N1534
  );


  not
  NOT1_439
  (
    N1593,
    N1537
  );


  nand
  NAND2_440
  (
    N1594,
    N1540,
    N1530
  );


  not
  NOT1_441
  (
    N1595,
    N1540
  );


  nand
  NAND2_442
  (
    N1596,
    N1567,
    N1568
  );


  buf
  BUFF1_443
  (
    N1600,
    N1517
  );


  buf
  BUFF1_444
  (
    N1603,
    N1517
  );


  buf
  BUFF1_445
  (
    N1606,
    N1522
  );


  buf
  BUFF1_446
  (
    N1609,
    N1522
  );


  buf
  BUFF1_447
  (
    N1612,
    N1514
  );


  buf
  BUFF1_448
  (
    N1615,
    N1514
  );


  buf
  BUFF1_449
  (
    N1620,
    N1557
  );


  buf
  BUFF1_450
  (
    N1623,
    N1554
  );


  not
  NOT1_451
  (
    N1635,
    N1571
  );


  nand
  NAND2_452
  (
    N1636,
    N1478,
    N1595
  );


  nand
  NAND2_453
  (
    N1638,
    N1576,
    N1569
  );


  not
  NOT1_454
  (
    N1639,
    N1576
  );


  buf
  BUFF1_455
  (
    N1640,
    N1561
  );


  buf
  BUFF1_456
  (
    N1643,
    N1561
  );


  buf
  BUFF1_457
  (
    N1647,
    N1546
  );


  buf
  BUFF1_458
  (
    N1651,
    N1546
  );


  buf
  BUFF1_459
  (
    N1658,
    N1554
  );


  buf
  BUFF1_460
  (
    N1661,
    N1557
  );


  buf
  BUFF1_461
  (
    N1664,
    N1557
  );


  nand
  NAND2_462
  (
    N1671,
    N1596,
    N893
  );


  not
  NOT1_463
  (
    N1672,
    N1596
  );


  not
  NOT1_464
  (
    N1675,
    N1600
  );


  not
  NOT1_465
  (
    N1677,
    N1603
  );


  nand
  NAND2_466
  (
    N1678,
    N1606,
    N1217
  );


  not
  NOT1_467
  (
    N1679,
    N1606
  );


  nand
  NAND2_468
  (
    N1680,
    N1609,
    N1219
  );


  not
  NOT1_469
  (
    N1681,
    N1609
  );


  not
  NOT1_470
  (
    N1682,
    N1612
  );


  not
  NOT1_471
  (
    N1683,
    N1615
  );


  nand
  NAND2_472
  (
    N1685,
    N1594,
    N1636
  );


  nand
  NAND2_473
  (
    N1688,
    N1510,
    N1639
  );


  buf
  BUFF1_474
  (
    N1697,
    N1588
  );


  buf
  BUFF1_475
  (
    N1701,
    N1588
  );


  nand
  NAND2_476
  (
    N1706,
    N643,
    N1672
  );


  not
  NOT1_477
  (
    N1707,
    N1643
  );


  nand
  NAND2_478
  (
    N1708,
    N1647,
    N1675
  );


  not
  NOT1_479
  (
    N1709,
    N1647
  );


  nand
  NAND2_480
  (
    N1710,
    N1651,
    N1677
  );


  not
  NOT1_481
  (
    N1711,
    N1651
  );


  nand
  NAND2_482
  (
    N1712,
    N1028,
    N1679
  );


  nand
  NAND2_483
  (
    N1713,
    N1031,
    N1681
  );


  buf
  BUFF1_484
  (
    N1714,
    N1620
  );


  buf
  BUFF1_485
  (
    N1717,
    N1620
  );


  nand
  NAND2_486
  (
    N1720,
    N1658,
    N1593
  );


  not
  NOT1_487
  (
    N1721,
    N1658
  );


  nand
  NAND2_488
  (
    N1723,
    N1638,
    N1688
  );


  not
  NOT1_489
  (
    N1727,
    N1661
  );


  not
  NOT1_490
  (
    N1728,
    N1640
  );


  not
  NOT1_491
  (
    N1730,
    N1664
  );


  buf
  BUFF1_492
  (
    N1731,
    N1623
  );


  buf
  BUFF1_493
  (
    N1734,
    N1623
  );


  nand
  NAND2_494
  (
    N1740,
    N1685,
    N1528
  );


  not
  NOT1_495
  (
    N1741,
    N1685
  );


  nand
  NAND2_496
  (
    N1742,
    N1671,
    N1706
  );


  nand
  NAND2_497
  (
    N1746,
    N1600,
    N1709
  );


  nand
  NAND2_498
  (
    N1747,
    N1603,
    N1711
  );


  nand
  NAND2_499
  (
    N1748,
    N1678,
    N1712
  );


  nand
  NAND2_500
  (
    N1751,
    N1680,
    N1713
  );


  nand
  NAND2_501
  (
    N1759,
    N1537,
    N1721
  );


  not
  NOT1_502
  (
    N1761,
    N1697
  );


  nand
  NAND2_503
  (
    N1762,
    N1697,
    N1727
  );


  not
  NOT1_504
  (
    N1763,
    N1701
  );


  nand
  NAND2_505
  (
    N1764,
    N1701,
    N1730
  );


  not
  NOT1_506
  (
    N1768,
    N1717
  );


  nand
  NAND2_507
  (
    N1769,
    N1472,
    N1741
  );


  nand
  NAND2_508
  (
    N1772,
    N1723,
    N1413
  );


  not
  NOT1_509
  (
    N1773,
    N1723
  );


  nand
  NAND2_510
  (
    N1774,
    N1708,
    N1746
  );


  nand
  NAND2_511
  (
    N1777,
    N1710,
    N1747
  );


  not
  NOT1_512
  (
    N1783,
    N1731
  );


  nand
  NAND2_513
  (
    N1784,
    N1731,
    N1682
  );


  not
  NOT1_514
  (
    N1785,
    N1714
  );


  not
  NOT1_515
  (
    N1786,
    N1734
  );


  nand
  NAND2_516
  (
    N1787,
    N1734,
    N1683
  );


  nand
  NAND2_517
  (
    N1788,
    N1720,
    N1759
  );


  nand
  NAND2_518
  (
    N1791,
    N1661,
    N1761
  );


  nand
  NAND2_519
  (
    N1792,
    N1664,
    N1763
  );


  nand
  NAND2_520
  (
    N1795,
    N1751,
    N1155
  );


  not
  NOT1_521
  (
    N1796,
    N1751
  );


  nand
  NAND2_522
  (
    N1798,
    N1740,
    N1769
  );


  nand
  NAND2_523
  (
    N1801,
    N1334,
    N1773
  );


  nand
  NAND2_524
  (
    N1802,
    N1742,
    N290
  );


  not
  NOT1_525
  (
    N1807,
    N1748
  );


  nand
  NAND2_526
  (
    N1808,
    N1748,
    N1218
  );


  nand
  NAND2_527
  (
    N1809,
    N1612,
    N1783
  );


  nand
  NAND2_528
  (
    N1810,
    N1615,
    N1786
  );


  nand
  NAND2_529
  (
    N1812,
    N1791,
    N1762
  );


  nand
  NAND2_530
  (
    N1815,
    N1792,
    N1764
  );


  buf
  BUFF1_531
  (
    N1818,
    N1742
  );


  nand
  NAND2_532
  (
    N1821,
    N1777,
    N1490
  );


  not
  NOT1_533
  (
    N1822,
    N1777
  );


  nand
  NAND2_534
  (
    N1823,
    N1774,
    N1491
  );


  not
  NOT1_535
  (
    N1824,
    N1774
  );


  nand
  NAND2_536
  (
    N1825,
    N962,
    N1796
  );


  nand
  NAND2_537
  (
    N1826,
    N1788,
    N1409
  );


  not
  NOT1_538
  (
    N1827,
    N1788
  );


  nand
  NAND2_539
  (
    N1830,
    N1772,
    N1801
  );


  nand
  NAND2_540
  (
    N1837,
    N959,
    N1807
  );


  nand
  NAND2_541
  (
    N1838,
    N1809,
    N1784
  );


  nand
  NAND2_542
  (
    N1841,
    N1810,
    N1787
  );


  nand
  NAND2_543
  (
    N1848,
    N1419,
    N1822
  );


  nand
  NAND2_544
  (
    N1849,
    N1416,
    N1824
  );


  nand
  NAND2_545
  (
    N1850,
    N1795,
    N1825
  );


  nand
  NAND2_546
  (
    N1852,
    N1319,
    N1827
  );


  nand
  NAND2_547
  (
    N1855,
    N1815,
    N1707
  );


  not
  NOT1_548
  (
    N1856,
    N1815
  );


  not
  NOT1_549
  (
    N1857,
    N1818
  );


  nand
  NAND2_550
  (
    N1858,
    N1798,
    N290
  );


  not
  NOT1_551
  (
    N1864,
    N1812
  );


  nand
  NAND2_552
  (
    N1865,
    N1812,
    N1728
  );


  buf
  BUFF1_553
  (
    N1866,
    N1798
  );


  buf
  BUFF1_554
  (
    N1869,
    N1802
  );


  buf
  BUFF1_555
  (
    N1872,
    N1802
  );


  nand
  NAND2_556
  (
    N1875,
    N1808,
    N1837
  );


  nand
  NAND2_557
  (
    N1878,
    N1821,
    N1848
  );


  nand
  NAND2_558
  (
    N1879,
    N1823,
    N1849
  );


  nand
  NAND2_559
  (
    N1882,
    N1841,
    N1768
  );


  not
  NOT1_560
  (
    N1883,
    N1841
  );


  nand
  NAND2_561
  (
    N1884,
    N1826,
    N1852
  );


  nand
  NAND2_562
  (
    N1885,
    N1643,
    N1856
  );


  nand
  NAND2_563
  (
    N1889,
    N1830,
    N290
  );


  not
  NOT1_564
  (
    N1895,
    N1838
  );


  nand
  NAND2_565
  (
    N1896,
    N1838,
    N1785
  );


  nand
  NAND2_566
  (
    N1897,
    N1640,
    N1864
  );


  not
  NOT1_567
  (
    N1898,
    N1850
  );


  buf
  BUFF1_568
  (
    N1902,
    N1830
  );


  not
  NOT1_569
  (
    N1910,
    N1878
  );


  nand
  NAND2_570
  (
    N1911,
    N1717,
    N1883
  );


  not
  NOT1_571
  (
    N1912,
    N1884
  );


  nand
  NAND2_572
  (
    N1913,
    N1855,
    N1885
  );


  not
  NOT1_573
  (
    N1915,
    N1866
  );


  nand
  NAND2_574
  (
    N1919,
    N1872,
    N919
  );


  not
  NOT1_575
  (
    N1920,
    N1872
  );


  nand
  NAND2_576
  (
    N1921,
    N1869,
    N920
  );


  not
  NOT1_577
  (
    N1922,
    N1869
  );


  not
  NOT1_578
  (
    N1923,
    N1875
  );


  nand
  NAND2_579
  (
    N1924,
    N1714,
    N1895
  );


  buf
  BUFF1_580
  (
    N1927,
    N1858
  );


  buf
  BUFF1_581
  (
    N1930,
    N1858
  );


  nand
  NAND2_582
  (
    N1933,
    N1865,
    N1897
  );


  nand
  NAND2_583
  (
    N1936,
    N1882,
    N1911
  );


  not
  NOT1_584
  (
    N1937,
    N1898
  );


  not
  NOT1_585
  (
    N1938,
    N1902
  );


  nand
  NAND2_586
  (
    N1941,
    N679,
    N1920
  );


  nand
  NAND2_587
  (
    N1942,
    N676,
    N1922
  );


  buf
  BUFF1_588
  (
    N1944,
    N1879
  );


  not
  NOT1_589
  (
    N1947,
    N1913
  );


  buf
  BUFF1_590
  (
    N1950,
    N1889
  );


  buf
  BUFF1_591
  (
    N1953,
    N1889
  );


  buf
  BUFF1_592
  (
    N1958,
    N1879
  );


  nand
  NAND2_593
  (
    N1961,
    N1896,
    N1924
  );


  and
  AND2_594
  (
    N1965,
    N1910,
    N601
  );


  and
  AND2_595
  (
    N1968,
    N602,
    N1912
  );


  nand
  NAND2_596
  (
    N1975,
    N1930,
    N917
  );


  not
  NOT1_597
  (
    N1976,
    N1930
  );


  nand
  NAND2_598
  (
    N1977,
    N1927,
    N918
  );


  not
  NOT1_599
  (
    N1978,
    N1927
  );


  nand
  NAND2_600
  (
    N1979,
    N1919,
    N1941
  );


  nand
  NAND2_601
  (
    N1980,
    N1921,
    N1942
  );


  not
  NOT1_602
  (
    N1985,
    N1933
  );


  not
  NOT1_603
  (
    N1987,
    N1936
  );


  not
  NOT1_604
  (
    N1999,
    N1944
  );


  nand
  NAND2_605
  (
    N2000,
    N1944,
    N1937
  );


  not
  NOT1_606
  (
    N2002,
    N1947
  );


  nand
  NAND2_607
  (
    N2003,
    N1947,
    N1499
  );


  nand
  NAND2_608
  (
    N2004,
    N1953,
    N1350
  );


  not
  NOT1_609
  (
    N2005,
    N1953
  );


  nand
  NAND2_610
  (
    N2006,
    N1950,
    N1351
  );


  not
  NOT1_611
  (
    N2007,
    N1950
  );


  nand
  NAND2_612
  (
    N2008,
    N673,
    N1976
  );


  nand
  NAND2_613
  (
    N2009,
    N670,
    N1978
  );


  not
  NOT1_614
  (
    N2012,
    N1979
  );


  not
  NOT1_615
  (
    N2013,
    N1958
  );


  nand
  NAND2_616
  (
    N2014,
    N1958,
    N1923
  );


  not
  NOT1_617
  (
    N2015,
    N1961
  );


  nand
  NAND2_618
  (
    N2016,
    N1961,
    N1635
  );


  not
  NOT1_619
  (
    N2018,
    N1965
  );


  not
  NOT1_620
  (
    N2019,
    N1968
  );


  nand
  NAND2_621
  (
    N2020,
    N1898,
    N1999
  );


  not
  NOT1_622
  (
    N2021,
    N1987
  );


  nand
  NAND2_623
  (
    N2022,
    N1987,
    N1591
  );


  nand
  NAND2_624
  (
    N2023,
    N1440,
    N2002
  );


  nand
  NAND2_625
  (
    N2024,
    N1261,
    N2005
  );


  nand
  NAND2_626
  (
    N2025,
    N1258,
    N2007
  );


  nand
  NAND2_627
  (
    N2026,
    N1975,
    N2008
  );


  nand
  NAND2_628
  (
    N2027,
    N1977,
    N2009
  );


  not
  NOT1_629
  (
    N2030,
    N1980
  );


  buf
  BUFF1_630
  (
    N2033,
    N1980
  );


  nand
  NAND2_631
  (
    N2036,
    N1875,
    N2013
  );


  nand
  NAND2_632
  (
    N2037,
    N1571,
    N2015
  );


  nand
  NAND2_633
  (
    N2038,
    N2020,
    N2000
  );


  nand
  NAND2_634
  (
    N2039,
    N1534,
    N2021
  );


  nand
  NAND2_635
  (
    N2040,
    N2023,
    N2003
  );


  nand
  NAND2_636
  (
    N2041,
    N2004,
    N2024
  );


  nand
  NAND2_637
  (
    N2042,
    N2006,
    N2025
  );


  not
  NOT1_638
  (
    N2047,
    N2026
  );


  nand
  NAND2_639
  (
    N2052,
    N2036,
    N2014
  );


  nand
  NAND2_640
  (
    N2055,
    N2037,
    N2016
  );


  not
  NOT1_641
  (
    N2060,
    N2038
  );


  nand
  NAND2_642
  (
    N2061,
    N2039,
    N2022
  );


  nand
  NAND2_643
  (
    N2062,
    N2040,
    N290
  );


  not
  NOT1_644
  (
    N2067,
    N2041
  );


  not
  NOT1_645
  (
    N2068,
    N2027
  );


  buf
  BUFF1_646
  (
    N2071,
    N2027
  );


  not
  NOT1_647
  (
    N2076,
    N2052
  );


  not
  NOT1_648
  (
    N2077,
    N2055
  );


  nand
  NAND2_649
  (
    N2078,
    N2060,
    N290
  );


  nand
  NAND2_650
  (
    N2081,
    N2061,
    N290
  );


  not
  NOT1_651
  (
    N2086,
    N2042
  );


  buf
  BUFF1_652
  (
    N2089,
    N2042
  );


  and
  AND2_653
  (
    N2104,
    N2030,
    N2068
  );


  and
  AND2_654
  (
    N2119,
    N2033,
    N2068
  );


  and
  AND2_655
  (
    N2129,
    N2030,
    N2071
  );


  and
  AND2_656
  (
    N2143,
    N2033,
    N2071
  );


  buf
  BUFF1_657
  (
    N2148,
    N2062
  );


  buf
  BUFF1_658
  (
    N2151,
    N2062
  );


  buf
  BUFF1_659
  (
    N2196,
    N2078
  );


  buf
  BUFF1_660
  (
    N2199,
    N2078
  );


  buf
  BUFF1_661
  (
    N2202,
    N2081
  );


  buf
  BUFF1_662
  (
    N2205,
    N2081
  );


  nand
  NAND2_663
  (
    N2214,
    N2151,
    N915
  );


  not
  NOT1_664
  (
    N2215,
    N2151
  );


  nand
  NAND2_665
  (
    N2216,
    N2148,
    N916
  );


  not
  NOT1_666
  (
    N2217,
    N2148
  );


  nand
  NAND2_667
  (
    N2222,
    N2199,
    N1348
  );


  not
  NOT1_668
  (
    N2223,
    N2199
  );


  nand
  NAND2_669
  (
    N2224,
    N2196,
    N1349
  );


  not
  NOT1_670
  (
    N2225,
    N2196
  );


  nand
  NAND2_671
  (
    N2226,
    N2205,
    N913
  );


  not
  NOT1_672
  (
    N2227,
    N2205
  );


  nand
  NAND2_673
  (
    N2228,
    N2202,
    N914
  );


  not
  NOT1_674
  (
    N2229,
    N2202
  );


  nand
  NAND2_675
  (
    N2230,
    N667,
    N2215
  );


  nand
  NAND2_676
  (
    N2231,
    N664,
    N2217
  );


  nand
  NAND2_677
  (
    N2232,
    N1255,
    N2223
  );


  nand
  NAND2_678
  (
    N2233,
    N1252,
    N2225
  );


  nand
  NAND2_679
  (
    N2234,
    N661,
    N2227
  );


  nand
  NAND2_680
  (
    N2235,
    N658,
    N2229
  );


  nand
  NAND2_681
  (
    N2236,
    N2214,
    N2230
  );


  nand
  NAND2_682
  (
    N2237,
    N2216,
    N2231
  );


  nand
  NAND2_683
  (
    N2240,
    N2222,
    N2232
  );


  nand
  NAND2_684
  (
    N2241,
    N2224,
    N2233
  );


  nand
  NAND2_685
  (
    N2244,
    N2226,
    N2234
  );


  nand
  NAND2_686
  (
    N2245,
    N2228,
    N2235
  );


  not
  NOT1_687
  (
    N2250,
    N2236
  );


  not
  NOT1_688
  (
    N2253,
    N2240
  );


  not
  NOT1_689
  (
    N2256,
    N2244
  );


  not
  NOT1_690
  (
    N2257,
    N2237
  );


  buf
  BUFF1_691
  (
    N2260,
    N2237
  );


  not
  NOT1_692
  (
    N2263,
    N2241
  );


  and
  AND2_693
  (
    N2266,
    N1164,
    N2241
  );


  not
  NOT1_694
  (
    N2269,
    N2245
  );


  and
  AND2_695
  (
    N2272,
    N1168,
    N2245
  );


  nand
  NAND8_696
  (
    N2279,
    N2067,
    N2012,
    N2047,
    N2250,
    N899,
    N2256,
    N2253,
    N903
  );


  buf
  BUFF1_697
  (
    N2286,
    N2266
  );


  buf
  BUFF1_698
  (
    N2297,
    N2266
  );


  buf
  BUFF1_699
  (
    N2315,
    N2272
  );


  buf
  BUFF1_700
  (
    N2326,
    N2272
  );


  and
  AND2_701
  (
    N2340,
    N2086,
    N2257
  );


  and
  AND2_702
  (
    N2353,
    N2089,
    N2257
  );


  and
  AND2_703
  (
    N2361,
    N2086,
    N2260
  );


  and
  AND2_704
  (
    N2375,
    N2089,
    N2260
  );


  and
  AND4_705
  (
    N2384,
    N338,
    N2279,
    N313,
    N313
  );


  and
  AND2_706
  (
    N2385,
    N1163,
    N2263
  );


  and
  AND2_707
  (
    N2386,
    N1164,
    N2263
  );


  and
  AND2_708
  (
    N2426,
    N1167,
    N2269
  );


  and
  AND2_709
  (
    N2427,
    N1168,
    N2269
  );


  nand
  NAND5_710
  (
    N2537,
    N2286,
    N2315,
    N2361,
    N2104,
    N1171
  );


  nand
  NAND5_711
  (
    N2540,
    N2286,
    N2315,
    N2340,
    N2129,
    N1171
  );


  nand
  NAND5_712
  (
    N2543,
    N2286,
    N2315,
    N2340,
    N2119,
    N1171
  );


  nand
  NAND5_713
  (
    N2546,
    N2286,
    N2315,
    N2353,
    N2104,
    N1171
  );


  nand
  NAND5_714
  (
    N2549,
    N2297,
    N2315,
    N2375,
    N2119,
    N1188
  );


  nand
  NAND5_715
  (
    N2552,
    N2297,
    N2326,
    N2361,
    N2143,
    N1188
  );


  nand
  NAND5_716
  (
    N2555,
    N2297,
    N2326,
    N2375,
    N2129,
    N1188
  );


  and
  AND5_717
  (
    N2558,
    N2286,
    N2315,
    N2361,
    N2104,
    N1171
  );


  and
  AND5_718
  (
    N2561,
    N2286,
    N2315,
    N2340,
    N2129,
    N1171
  );


  and
  AND5_719
  (
    N2564,
    N2286,
    N2315,
    N2340,
    N2119,
    N1171
  );


  and
  AND5_720
  (
    N2567,
    N2286,
    N2315,
    N2353,
    N2104,
    N1171
  );


  and
  AND5_721
  (
    N2570,
    N2297,
    N2315,
    N2375,
    N2119,
    N1188
  );


  and
  AND5_722
  (
    N2573,
    N2297,
    N2326,
    N2361,
    N2143,
    N1188
  );


  and
  AND5_723
  (
    N2576,
    N2297,
    N2326,
    N2375,
    N2129,
    N1188
  );


  nand
  NAND5_724
  (
    N2594,
    N2286,
    N2427,
    N2361,
    N2129,
    N1171
  );


  nand
  NAND5_725
  (
    N2597,
    N2297,
    N2427,
    N2361,
    N2119,
    N1171
  );


  nand
  NAND5_726
  (
    N2600,
    N2297,
    N2427,
    N2375,
    N2104,
    N1171
  );


  nand
  NAND5_727
  (
    N2603,
    N2297,
    N2427,
    N2340,
    N2143,
    N1171
  );


  nand
  NAND5_728
  (
    N2606,
    N2297,
    N2427,
    N2353,
    N2129,
    N1188
  );


  nand
  NAND5_729
  (
    N2611,
    N2386,
    N2326,
    N2361,
    N2129,
    N1188
  );


  nand
  NAND5_730
  (
    N2614,
    N2386,
    N2326,
    N2361,
    N2119,
    N1188
  );


  nand
  NAND5_731
  (
    N2617,
    N2386,
    N2326,
    N2375,
    N2104,
    N1188
  );


  nand
  NAND5_732
  (
    N2620,
    N2386,
    N2326,
    N2353,
    N2129,
    N1188
  );


  nand
  NAND5_733
  (
    N2627,
    N2297,
    N2427,
    N2340,
    N2104,
    N926
  );


  nand
  NAND5_734
  (
    N2628,
    N2386,
    N2326,
    N2340,
    N2104,
    N926
  );


  nand
  NAND5_735
  (
    N2629,
    N2386,
    N2427,
    N2361,
    N2104,
    N926
  );


  nand
  NAND5_736
  (
    N2630,
    N2386,
    N2427,
    N2340,
    N2129,
    N926
  );


  nand
  NAND5_737
  (
    N2631,
    N2386,
    N2427,
    N2340,
    N2119,
    N926
  );


  nand
  NAND5_738
  (
    N2632,
    N2386,
    N2427,
    N2353,
    N2104,
    N926
  );


  nand
  NAND5_739
  (
    N2633,
    N2386,
    N2426,
    N2340,
    N2104,
    N926
  );


  nand
  NAND5_740
  (
    N2634,
    N2385,
    N2427,
    N2340,
    N2104,
    N926
  );


  and
  AND5_741
  (
    N2639,
    N2286,
    N2427,
    N2361,
    N2129,
    N1171
  );


  and
  AND5_742
  (
    N2642,
    N2297,
    N2427,
    N2361,
    N2119,
    N1171
  );


  and
  AND5_743
  (
    N2645,
    N2297,
    N2427,
    N2375,
    N2104,
    N1171
  );


  and
  AND5_744
  (
    N2648,
    N2297,
    N2427,
    N2340,
    N2143,
    N1171
  );


  and
  AND5_745
  (
    N2651,
    N2297,
    N2427,
    N2353,
    N2129,
    N1188
  );


  and
  AND5_746
  (
    N2655,
    N2386,
    N2326,
    N2361,
    N2129,
    N1188
  );


  and
  AND5_747
  (
    N2658,
    N2386,
    N2326,
    N2361,
    N2119,
    N1188
  );


  and
  AND5_748
  (
    N2661,
    N2386,
    N2326,
    N2375,
    N2104,
    N1188
  );


  and
  AND5_749
  (
    N2664,
    N2386,
    N2326,
    N2353,
    N2129,
    N1188
  );


  nand
  NAND2_750
  (
    N2669,
    N2558,
    N534
  );


  not
  NOT1_751
  (
    N2670,
    N2558
  );


  nand
  NAND2_752
  (
    N2671,
    N2561,
    N535
  );


  not
  NOT1_753
  (
    N2672,
    N2561
  );


  nand
  NAND2_754
  (
    N2673,
    N2564,
    N536
  );


  not
  NOT1_755
  (
    N2674,
    N2564
  );


  nand
  NAND2_756
  (
    N2675,
    N2567,
    N537
  );


  not
  NOT1_757
  (
    N2676,
    N2567
  );


  nand
  NAND2_758
  (
    N2682,
    N2570,
    N543
  );


  not
  NOT1_759
  (
    N2683,
    N2570
  );


  nand
  NAND2_760
  (
    N2688,
    N2573,
    N548
  );


  not
  NOT1_761
  (
    N2689,
    N2573
  );


  nand
  NAND2_762
  (
    N2690,
    N2576,
    N549
  );


  not
  NOT1_763
  (
    N2691,
    N2576
  );


  and
  AND8_764
  (
    N2710,
    N2627,
    N2628,
    N2629,
    N2630,
    N2631,
    N2632,
    N2633,
    N2634
  );


  nand
  NAND2_765
  (
    N2720,
    N343,
    N2670
  );


  nand
  NAND2_766
  (
    N2721,
    N346,
    N2672
  );


  nand
  NAND2_767
  (
    N2722,
    N349,
    N2674
  );


  nand
  NAND2_768
  (
    N2723,
    N352,
    N2676
  );


  nand
  NAND2_769
  (
    N2724,
    N2639,
    N538
  );


  not
  NOT1_770
  (
    N2725,
    N2639
  );


  nand
  NAND2_771
  (
    N2726,
    N2642,
    N539
  );


  not
  NOT1_772
  (
    N2727,
    N2642
  );


  nand
  NAND2_773
  (
    N2728,
    N2645,
    N540
  );


  not
  NOT1_774
  (
    N2729,
    N2645
  );


  nand
  NAND2_775
  (
    N2730,
    N2648,
    N541
  );


  not
  NOT1_776
  (
    N2731,
    N2648
  );


  nand
  NAND2_777
  (
    N2732,
    N2651,
    N542
  );


  not
  NOT1_778
  (
    N2733,
    N2651
  );


  nand
  NAND2_779
  (
    N2734,
    N370,
    N2683
  );


  nand
  NAND2_780
  (
    N2735,
    N2655,
    N544
  );


  not
  NOT1_781
  (
    N2736,
    N2655
  );


  nand
  NAND2_782
  (
    N2737,
    N2658,
    N545
  );


  not
  NOT1_783
  (
    N2738,
    N2658
  );


  nand
  NAND2_784
  (
    N2739,
    N2661,
    N546
  );


  not
  NOT1_785
  (
    N2740,
    N2661
  );


  nand
  NAND2_786
  (
    N2741,
    N2664,
    N547
  );


  not
  NOT1_787
  (
    N2742,
    N2664
  );


  nand
  NAND2_788
  (
    N2743,
    N385,
    N2689
  );


  nand
  NAND2_789
  (
    N2744,
    N388,
    N2691
  );


  nand
  NAND8_790
  (
    N2745,
    N2537,
    N2540,
    N2543,
    N2546,
    N2594,
    N2597,
    N2600,
    N2603
  );


  nand
  NAND8_791
  (
    N2746,
    N2606,
    N2549,
    N2611,
    N2614,
    N2617,
    N2620,
    N2552,
    N2555
  );


  and
  AND8_792
  (
    N2747,
    N2537,
    N2540,
    N2543,
    N2546,
    N2594,
    N2597,
    N2600,
    N2603
  );


  and
  AND8_793
  (
    N2750,
    N2606,
    N2549,
    N2611,
    N2614,
    N2617,
    N2620,
    N2552,
    N2555
  );


  nand
  NAND2_794
  (
    N2753,
    N2669,
    N2720
  );


  nand
  NAND2_795
  (
    N2754,
    N2671,
    N2721
  );


  nand
  NAND2_796
  (
    N2755,
    N2673,
    N2722
  );


  nand
  NAND2_797
  (
    N2756,
    N2675,
    N2723
  );


  nand
  NAND2_798
  (
    N2757,
    N355,
    N2725
  );


  nand
  NAND2_799
  (
    N2758,
    N358,
    N2727
  );


  nand
  NAND2_800
  (
    N2759,
    N361,
    N2729
  );


  nand
  NAND2_801
  (
    N2760,
    N364,
    N2731
  );


  nand
  NAND2_802
  (
    N2761,
    N367,
    N2733
  );


  nand
  NAND2_803
  (
    N2762,
    N2682,
    N2734
  );


  nand
  NAND2_804
  (
    N2763,
    N373,
    N2736
  );


  nand
  NAND2_805
  (
    N2764,
    N376,
    N2738
  );


  nand
  NAND2_806
  (
    N2765,
    N379,
    N2740
  );


  nand
  NAND2_807
  (
    N2766,
    N382,
    N2742
  );


  nand
  NAND2_808
  (
    N2767,
    N2688,
    N2743
  );


  nand
  NAND2_809
  (
    N2768,
    N2690,
    N2744
  );


  and
  AND2_810
  (
    N2773,
    N2745,
    N275
  );


  and
  AND2_811
  (
    N2776,
    N2746,
    N276
  );


  nand
  NAND2_812
  (
    N2779,
    N2724,
    N2757
  );


  nand
  NAND2_813
  (
    N2780,
    N2726,
    N2758
  );


  nand
  NAND2_814
  (
    N2781,
    N2728,
    N2759
  );


  nand
  NAND2_815
  (
    N2782,
    N2730,
    N2760
  );


  nand
  NAND2_816
  (
    N2783,
    N2732,
    N2761
  );


  nand
  NAND2_817
  (
    N2784,
    N2735,
    N2763
  );


  nand
  NAND2_818
  (
    N2785,
    N2737,
    N2764
  );


  nand
  NAND2_819
  (
    N2786,
    N2739,
    N2765
  );


  nand
  NAND2_820
  (
    N2787,
    N2741,
    N2766
  );


  and
  AND3_821
  (
    N2788,
    N2747,
    N2750,
    N2710
  );


  nand
  NAND2_822
  (
    N2789,
    N2747,
    N2750
  );


  and
  AND4_823
  (
    N2800,
    N338,
    N2279,
    N99,
    N2788
  );


  nand
  NAND2_824
  (
    N2807,
    N2773,
    N2018
  );


  not
  NOT1_825
  (
    N2808,
    N2773
  );


  nand
  NAND2_826
  (
    N2809,
    N2776,
    N2019
  );


  not
  NOT1_827
  (
    N2810,
    N2776
  );


  nor
  NOR2_828
  (
    N2811,
    N2384,
    N2800
  );


  and
  AND3_829
  (
    N2812,
    N897,
    N283,
    N2789
  );


  and
  AND3_830
  (
    N2815,
    N76,
    N283,
    N2789
  );


  and
  AND3_831
  (
    N2818,
    N82,
    N283,
    N2789
  );


  and
  AND3_832
  (
    N2821,
    N85,
    N283,
    N2789
  );


  and
  AND3_833
  (
    N2824,
    N898,
    N283,
    N2789
  );


  nand
  NAND2_834
  (
    N2827,
    N1965,
    N2808
  );


  nand
  NAND2_835
  (
    N2828,
    N1968,
    N2810
  );


  and
  AND3_836
  (
    N2829,
    N79,
    N283,
    N2789
  );


  nand
  NAND2_837
  (
    N2843,
    N2807,
    N2827
  );


  nand
  NAND2_838
  (
    N2846,
    N2809,
    N2828
  );


  nand
  NAND2_839
  (
    N2850,
    N2812,
    N2076
  );


  nand
  NAND2_840
  (
    N2851,
    N2815,
    N2077
  );


  nand
  NAND2_841
  (
    N2852,
    N2818,
    N1915
  );


  nand
  NAND2_842
  (
    N2853,
    N2821,
    N1857
  );


  nand
  NAND2_843
  (
    N2854,
    N2824,
    N1938
  );


  not
  NOT1_844
  (
    N2857,
    N2812
  );


  not
  NOT1_845
  (
    N2858,
    N2815
  );


  not
  NOT1_846
  (
    N2859,
    N2818
  );


  not
  NOT1_847
  (
    N2860,
    N2821
  );


  not
  NOT1_848
  (
    N2861,
    N2824
  );


  not
  NOT1_849
  (
    N2862,
    N2829
  );


  nand
  NAND2_850
  (
    N2863,
    N2829,
    N1985
  );


  nand
  NAND2_851
  (
    N2866,
    N2052,
    N2857
  );


  nand
  NAND2_852
  (
    N2867,
    N2055,
    N2858
  );


  nand
  NAND2_853
  (
    N2868,
    N1866,
    N2859
  );


  nand
  NAND2_854
  (
    N2869,
    N1818,
    N2860
  );


  nand
  NAND2_855
  (
    N2870,
    N1902,
    N2861
  );


  nand
  NAND2_856
  (
    N2871,
    N2843,
    N886
  );


  not
  NOT1_857
  (
    N2872,
    N2843
  );


  nand
  NAND2_858
  (
    N2873,
    N2846,
    N887
  );


  not
  NOT1_859
  (
    N2874,
    N2846
  );


  nand
  NAND2_860
  (
    N2875,
    N1933,
    N2862
  );


  nand
  NAND2_861
  (
    N2876,
    N2866,
    N2850
  );


  nand
  NAND2_862
  (
    N2877,
    N2867,
    N2851
  );


  nand
  NAND2_863
  (
    N2878,
    N2868,
    N2852
  );


  nand
  NAND2_864
  (
    N2879,
    N2869,
    N2853
  );


  nand
  NAND2_865
  (
    N2880,
    N2870,
    N2854
  );


  nand
  NAND2_866
  (
    N2881,
    N682,
    N2872
  );


  nand
  NAND2_867
  (
    N2882,
    N685,
    N2874
  );


  nand
  NAND2_868
  (
    N2883,
    N2875,
    N2863
  );


  and
  AND2_869
  (
    signal_from_circuit_0,
    N2876,
    N550
  );


  and
  AND2_870
  (
    N2887,
    N551,
    N2877
  );


  and
  AND2_871
  (
    N2888,
    N553,
    N2878
  );


  and
  AND2_872
  (
    N2889,
    N2879,
    N554
  );


  and
  AND2_873
  (
    N2890,
    N555,
    N2880
  );


  nand
  NAND2_874
  (
    N2891,
    N2871,
    N2881
  );


  nand
  NAND2_875
  (
    N2892,
    N2873,
    N2882
  );


  nand
  NAND2_876
  (
    N2895,
    N2883,
    N1461
  );


  not
  NOT1_877
  (
    N2896,
    N2883
  );


  nand
  NAND2_878
  (
    N2897,
    N1383,
    N2896
  );


  nand
  NAND2_879
  (
    N2898,
    N2895,
    N2897
  );


  and
  AND2_880
  (
    N2899,
    N2898,
    N552
  );


  xnor
  SIG_COMP_XOR_0_0
  (
    sig_comp_0_0,
    keyIn_0_0,
    N1
  );


  xnor
  SIG_COMP_XOR_0_1
  (
    sig_comp_0_1,
    keyIn_0_1,
    N4
  );


  xnor
  SIG_COMP_XOR_0_2
  (
    sig_comp_0_2,
    keyIn_0_2,
    N7
  );


  xnor
  SIG_COMP_XOR_0_3
  (
    sig_comp_0_3,
    keyIn_0_3,
    N10
  );


  xnor
  SIG_COMP_XOR_0_4
  (
    sig_comp_0_4,
    keyIn_0_4,
    N13
  );


  xnor
  SIG_COMP_XOR_0_5
  (
    sig_comp_0_5,
    keyIn_0_5,
    N16
  );


  xnor
  SIG_COMP_XOR_0_6
  (
    sig_comp_0_6,
    keyIn_0_6,
    N19
  );


  xnor
  SIG_COMP_XOR_0_7
  (
    sig_comp_0_7,
    keyIn_0_7,
    N22
  );


  and
  SIG_COMP_AND_0
  (
    sig_comp_and_0,
    sig_comp_0_0,
    sig_comp_0_1,
    sig_comp_0_2,
    sig_comp_0_3,
    sig_comp_0_4,
    sig_comp_0_5,
    sig_comp_0_6,
    sig_comp_0_7
  );


  xnor
  CONST_COMP_XOR_0_0
  (
    const_comp_xor_0_0,
    keyIn_0_0,
    0
  );


  xnor
  CONST_COMP_XOR_0_1
  (
    const_comp_xor_0_1,
    keyIn_0_1,
    0
  );


  xnor
  CONST_COMP_XOR_0_2
  (
    const_comp_xor_0_2,
    keyIn_0_2,
    0
  );


  xnor
  CONST_COMP_XOR_0_3
  (
    const_comp_xor_0_3,
    keyIn_0_3,
    0
  );


  xnor
  CONST_COMP_XOR_0_4
  (
    const_comp_xor_0_4,
    keyIn_0_4,
    0
  );


  xnor
  CONST_COMP_XOR_0_5
  (
    const_comp_xor_0_5,
    keyIn_0_5,
    0
  );


  xnor
  CONST_COMP_XOR_0_6
  (
    const_comp_xor_0_6,
    keyIn_0_6,
    0
  );


  xnor
  CONST_COMP_XOR_0_7
  (
    const_comp_xor_0_7,
    keyIn_0_7,
    0
  );


  and
  CONST_COMP_AND_0
  (
    const_comp_and_0,
    const_comp_xor_0_0,
    const_comp_xor_0_1,
    const_comp_xor_0_2,
    const_comp_xor_0_3,
    const_comp_xor_0_4,
    const_comp_xor_0_5,
    const_comp_xor_0_6,
    const_comp_xor_0_7
  );


  and
  MASK_AND_0
  (
    mask_and_0,
    sig_comp_and_0,
    const_comp_and_0
  );


  xor
  FLIP_IT_0
  (
    flipped_signal_1,
    mask_and_0,
    signal_from_circuit_0
  );


  xor
  MUX_CONTROL_XOR_1_0
  (
    mux_control_xor_1_0,
    keyIn_1_8,
    N25
  );


  xor
  MUX_CONTROL_XOR_1_1
  (
    mux_control_xor_1_1,
    keyIn_1_9,
    N28
  );


  not
  MUX_NOT_1_0
  (
    mux_not_1_0,
    mux_control_xor_1_0
  );


  and
  MUX_AND0_1_0
  (
    mux_and0_1_0,
    signal_from_circuit_0,
    mux_not_1_0
  );


  and
  MUX_AND1_1_0
  (
    mux_and1_1_0,
    flipped_signal_1,
    mux_control_xor_1_0
  );


  or
  MUX_OR_1_0
  (
    mux_output_0,
    mux_and0_1_0,
    mux_and1_1_0
  );


  not
  MUX_NOT_1_1
  (
    mux_not_1_1,
    mux_control_xor_1_1
  );


  and
  MUX_AND0_1_1
  (
    mux_and0_1_1,
    signal_from_circuit_0,
    mux_not_1_1
  );


  and
  MUX_AND1_1_1
  (
    mux_and1_1_1,
    mux_output_0,
    mux_control_xor_1_1
  );


  or
  MUX_OR_1_1
  (
    N2886,
    mux_and0_1_1,
    mux_and1_1_1
  );


endmodule

